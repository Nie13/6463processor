----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:10:08 12/02/2017 
-- Design Name: 
-- Module Name:    Counter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY Counter IS

PORT 
	(	input : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		output : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		clk : IN STD_LOGIC;
		clr : IN STD_LOGIC
	);

END Counter;

ARCHITECTURE Behavioral OF Counter IS

BEGIN

	PROCESS (clk, input) 
	BEGIN
		IF(clk'EVENT AND clk = '1') THEN
			IF (clr = '1') THEN
				output <= (OTHERS =>'0');
			ELSE		
				output <= input;
			END IF;
		END IF;	
	END PROCESS;

END Behavioral;